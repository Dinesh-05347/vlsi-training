module and_gate_p (output c,input a, b);
and andg(c,a,b);
endmodule